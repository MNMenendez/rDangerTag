----------------------------------------------------------------------------------
-- Company: 
-- Engineer: 
-- 
-- Create Date:    14:27:43 05/01/2023 
-- Design Name: 
-- Module Name:    POWER - POWER_FUNC 
-- Project Name: 
-- Target Devices: 
-- Tool versions: 
-- Description: 
--
-- Dependencies: 
--
-- Revision: 
-- Revision 0.01 - File Created
-- Additional Comments: 
--
----------------------------------------------------------------------------------
library IEEE;
use IEEE.STD_LOGIC_1164.ALL;

-- Uncomment the following library declaration if using
-- arithmetic functions with Signed or Unsigned values
--use IEEE.NUMERIC_STD.ALL;

-- Uncomment the following library declaration if instantiating
-- any Xilinx primitives in this code.
--library UNISIM;
--use UNISIM.VComponents.all;

entity POWER_MODULE is
    Port ( PWR : in  STD_LOGIC;
           PWR_STATE : out  STD_LOGIC);
end POWER_MODULE;

architecture POWER_FUNC of POWER_MODULE is

begin


end POWER_FUNC;

