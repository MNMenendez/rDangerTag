----------------------------------------------------------------------------------
-- Company: 
-- Engineer: 
-- 
-- Create Date:    09:38:38 05/02/2023 
-- Design Name: 
-- Module Name:    DUMMY_MODULE - Behavioral 
-- Project Name: 
-- Target Devices: 
-- Tool versions: 
-- Description: 
--
-- Dependencies: 
--
-- Revision: 
-- Revision 0.01 - File Created
-- Additional Comments: 
--
----------------------------------------------------------------------------------
library IEEE;
use IEEE.STD_LOGIC_1164.ALL;

-- Uncomment the following library declaration if using
-- arithmetic functions with Signed or Unsigned values
--use IEEE.NUMERIC_STD.ALL;

-- Uncomment the following library declaration if instantiating
-- any Xilinx primitives in this code.
--library UNISIM;
--use UNISIM.VComponents.all;

entity DUMMY_MODULE is
    Port ( TBD_I : in  STD_LOGIC;
           TBD_O : out  STD_LOGIC);
end DUMMY_MODULE;

architecture DUMMY_FUNC of DUMMY_MODULE is

begin


end DUMMY_FUNC;

